library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity window_table is
	port (
		address : in std_logic_vector(11 downto 0);-- table address
		window_val : out std_logic_vector(11 downto 0)-- table entry value
		);
end window_table;

architecture behavioral of window_table is
	type lut is array(0 to 4095) of std_logic_vector(11 downto 0);
		constant window_lut : lut := (
"000011011101","000011011101","000011011110","000011011110","000011011110","000011011111","000011011111","000011100000","000011100000","000011100001",
"000011100001","000011100001","000011100010","000011100010","000011100011","000011100011","000011100100","000011100100","000011100101","000011100101",
"000011100101","000011100110","000011100110","000011100111","000011100111","000011101000","000011101000","000011101001","000011101001","000011101001",
"000011101010","000011101010","000011101011","000011101011","000011101100","000011101100","000011101101","000011101101","000011101110","000011101110",
"000011101110","000011101111","000011101111","000011110000","000011110000","000011110001","000011110001","000011110010","000011110010","000011110011",
"000011110011","000011110100","000011110100","000011110100","000011110101","000011110101","000011110110","000011110110","000011110111","000011110111",
"000011111000","000011111000","000011111001","000011111001","000011111010","000011111010","000011111011","000011111011","000011111100","000011111100",
"000011111100","000011111101","000011111101","000011111110","000011111110","000011111111","000011111111","000100000000","000100000000","000100000001",
"000100000001","000100000010","000100000010","000100000011","000100000011","000100000100","000100000100","000100000101","000100000101","000100000110",
"000100000110","000100000111","000100000111","000100001000","000100001000","000100001001","000100001001","000100001010","000100001010","000100001011",
"000100001011","000100001100","000100001100","000100001101","000100001101","000100001110","000100001110","000100001111","000100001111","000100010000",
"000100010000","000100010001","000100010001","000100010010","000100010010","000100010011","000100010011","000100010100","000100010100","000100010101",
"000100010101","000100010110","000100010110","000100010111","000100010111","000100011000","000100011000","000100011001","000100011001","000100011010",
"000100011010","000100011011","000100011011","000100011100","000100011100","000100011101","000100011101","000100011110","000100011110","000100011111",
"000100011111","000100100000","000100100001","000100100001","000100100010","000100100010","000100100011","000100100011","000100100100","000100100100",
"000100100101","000100100101","000100100110","000100100110","000100100111","000100100111","000100101000","000100101000","000100101001","000100101010",
"000100101010","000100101011","000100101011","000100101100","000100101100","000100101101","000100101101","000100101110","000100101110","000100101111",
"000100110000","000100110000","000100110001","000100110001","000100110010","000100110010","000100110011","000100110011","000100110100","000100110100",
"000100110101","000100110110","000100110110","000100110111","000100110111","000100111000","000100111000","000100111001","000100111001","000100111010",
"000100111011","000100111011","000100111100","000100111100","000100111101","000100111101","000100111110","000100111110","000100111111","000101000000",
"000101000000","000101000001","000101000001","000101000010","000101000010","000101000011","000101000100","000101000100","000101000101","000101000101",
"000101000110","000101000110","000101000111","000101001000","000101001000","000101001001","000101001001","000101001010","000101001010","000101001011",
"000101001100","000101001100","000101001101","000101001101","000101001110","000101001111","000101001111","000101010000","000101010000","000101010001",
"000101010001","000101010010","000101010011","000101010011","000101010100","000101010100","000101010101","000101010110","000101010110","000101010111",
"000101010111","000101011000","000101011001","000101011001","000101011010","000101011010","000101011011","000101011011","000101011100","000101011101",
"000101011101","000101011110","000101011110","000101011111","000101100000","000101100000","000101100001","000101100001","000101100010","000101100011",
"000101100011","000101100100","000101100101","000101100101","000101100110","000101100110","000101100111","000101101000","000101101000","000101101001",
"000101101001","000101101010","000101101011","000101101011","000101101100","000101101100","000101101101","000101101110","000101101110","000101101111",
"000101110000","000101110000","000101110001","000101110001","000101110010","000101110011","000101110011","000101110100","000101110101","000101110101",
"000101110110","000101110110","000101110111","000101111000","000101111000","000101111001","000101111010","000101111010","000101111011","000101111100",
"000101111100","000101111101","000101111101","000101111110","000101111111","000101111111","000110000000","000110000001","000110000001","000110000010",
"000110000011","000110000011","000110000100","000110000100","000110000101","000110000110","000110000110","000110000111","000110001000","000110001000",
"000110001001","000110001010","000110001010","000110001011","000110001100","000110001100","000110001101","000110001110","000110001110","000110001111",
"000110001111","000110010000","000110010001","000110010001","000110010010","000110010011","000110010011","000110010100","000110010101","000110010101",
"000110010110","000110010111","000110010111","000110011000","000110011001","000110011001","000110011010","000110011011","000110011011","000110011100",
"000110011101","000110011101","000110011110","000110011111","000110011111","000110100000","000110100001","000110100001","000110100010","000110100011",
"000110100011","000110100100","000110100101","000110100101","000110100110","000110100111","000110101000","000110101000","000110101001","000110101010",
"000110101010","000110101011","000110101100","000110101100","000110101101","000110101110","000110101110","000110101111","000110110000","000110110000",
"000110110001","000110110010","000110110010","000110110011","000110110100","000110110101","000110110101","000110110110","000110110111","000110110111",
"000110111000","000110111001","000110111001","000110111010","000110111011","000110111100","000110111100","000110111101","000110111110","000110111110",
"000110111111","000111000000","000111000000","000111000001","000111000010","000111000011","000111000011","000111000100","000111000101","000111000101",
"000111000110","000111000111","000111001000","000111001000","000111001001","000111001010","000111001010","000111001011","000111001100","000111001101",
"000111001101","000111001110","000111001111","000111001111","000111010000","000111010001","000111010010","000111010010","000111010011","000111010100",
"000111010100","000111010101","000111010110","000111010111","000111010111","000111011000","000111011001","000111011010","000111011010","000111011011",
"000111011100","000111011100","000111011101","000111011110","000111011111","000111011111","000111100000","000111100001","000111100010","000111100010",
"000111100011","000111100100","000111100101","000111100101","000111100110","000111100111","000111100111","000111101000","000111101001","000111101010",
"000111101010","000111101011","000111101100","000111101101","000111101101","000111101110","000111101111","000111110000","000111110000","000111110001",
"000111110010","000111110011","000111110011","000111110100","000111110101","000111110110","000111110110","000111110111","000111111000","000111111001",
"000111111001","000111111010","000111111011","000111111100","000111111100","000111111101","000111111110","000111111111","001000000000","001000000000",
"001000000001","001000000010","001000000011","001000000011","001000000100","001000000101","001000000110","001000000110","001000000111","001000001000",
"001000001001","001000001001","001000001010","001000001011","001000001100","001000001101","001000001101","001000001110","001000001111","001000010000",
"001000010000","001000010001","001000010010","001000010011","001000010100","001000010100","001000010101","001000010110","001000010111","001000010111",
"001000011000","001000011001","001000011010","001000011011","001000011011","001000011100","001000011101","001000011110","001000011111","001000011111",
"001000100000","001000100001","001000100010","001000100010","001000100011","001000100100","001000100101","001000100110","001000100110","001000100111",
"001000101000","001000101001","001000101010","001000101010","001000101011","001000101100","001000101101","001000101110","001000101110","001000101111",
"001000110000","001000110001","001000110010","001000110010","001000110011","001000110100","001000110101","001000110110","001000110110","001000110111",
"001000111000","001000111001","001000111010","001000111010","001000111011","001000111100","001000111101","001000111110","001000111110","001000111111",
"001001000000","001001000001","001001000010","001001000011","001001000011","001001000100","001001000101","001001000110","001001000111","001001000111",
"001001001000","001001001001","001001001010","001001001011","001001001100","001001001100","001001001101","001001001110","001001001111","001001010000",
"001001010000","001001010001","001001010010","001001010011","001001010100","001001010101","001001010101","001001010110","001001010111","001001011000",
"001001011001","001001011010","001001011010","001001011011","001001011100","001001011101","001001011110","001001011111","001001011111","001001100000",
"001001100001","001001100010","001001100011","001001100100","001001100100","001001100101","001001100110","001001100111","001001101000","001001101001",
"001001101001","001001101010","001001101011","001001101100","001001101101","001001101110","001001101111","001001101111","001001110000","001001110001",
"001001110010","001001110011","001001110100","001001110100","001001110101","001001110110","001001110111","001001111000","001001111001","001001111010",
"001001111010","001001111011","001001111100","001001111101","001001111110","001001111111","001010000000","001010000000","001010000001","001010000010",
"001010000011","001010000100","001010000101","001010000110","001010000110","001010000111","001010001000","001010001001","001010001010","001010001011",
"001010001100","001010001100","001010001101","001010001110","001010001111","001010010000","001010010001","001010010010","001010010011","001010010011",
"001010010100","001010010101","001010010110","001010010111","001010011000","001010011001","001010011001","001010011010","001010011011","001010011100",
"001010011101","001010011110","001010011111","001010100000","001010100000","001010100001","001010100010","001010100011","001010100100","001010100101",
"001010100110","001010100111","001010100111","001010101000","001010101001","001010101010","001010101011","001010101100","001010101101","001010101110",
"001010101111","001010101111","001010110000","001010110001","001010110010","001010110011","001010110100","001010110101","001010110110","001010110110",
"001010110111","001010111000","001010111001","001010111010","001010111011","001010111100","001010111101","001010111110","001010111110","001010111111",
"001011000000","001011000001","001011000010","001011000011","001011000100","001011000101","001011000110","001011000111","001011000111","001011001000",
"001011001001","001011001010","001011001011","001011001100","001011001101","001011001110","001011001111","001011010000","001011010000","001011010001",
"001011010010","001011010011","001011010100","001011010101","001011010110","001011010111","001011011000","001011011001","001011011001","001011011010",
"001011011011","001011011100","001011011101","001011011110","001011011111","001011100000","001011100001","001011100010","001011100011","001011100011",
"001011100100","001011100101","001011100110","001011100111","001011101000","001011101001","001011101010","001011101011","001011101100","001011101101",
"001011101101","001011101110","001011101111","001011110000","001011110001","001011110010","001011110011","001011110100","001011110101","001011110110",
"001011110111","001011111000","001011111000","001011111001","001011111010","001011111011","001011111100","001011111101","001011111110","001011111111",
"001100000000","001100000001","001100000010","001100000011","001100000100","001100000100","001100000101","001100000110","001100000111","001100001000",
"001100001001","001100001010","001100001011","001100001100","001100001101","001100001110","001100001111","001100010000","001100010000","001100010001",
"001100010010","001100010011","001100010100","001100010101","001100010110","001100010111","001100011000","001100011001","001100011010","001100011011",
"001100011100","001100011101","001100011101","001100011110","001100011111","001100100000","001100100001","001100100010","001100100011","001100100100",
"001100100101","001100100110","001100100111","001100101000","001100101001","001100101010","001100101011","001100101100","001100101100","001100101101",
"001100101110","001100101111","001100110000","001100110001","001100110010","001100110011","001100110100","001100110101","001100110110","001100110111",
"001100111000","001100111001","001100111010","001100111011","001100111100","001100111100","001100111101","001100111110","001100111111","001101000000",
"001101000001","001101000010","001101000011","001101000100","001101000101","001101000110","001101000111","001101001000","001101001001","001101001010",
"001101001011","001101001100","001101001101","001101001101","001101001110","001101001111","001101010000","001101010001","001101010010","001101010011",
"001101010100","001101010101","001101010110","001101010111","001101011000","001101011001","001101011010","001101011011","001101011100","001101011101",
"001101011110","001101011111","001101100000","001101100000","001101100001","001101100010","001101100011","001101100100","001101100101","001101100110",
"001101100111","001101101000","001101101001","001101101010","001101101011","001101101100","001101101101","001101101110","001101101111","001101110000",
"001101110001","001101110010","001101110011","001101110100","001101110101","001101110110","001101110110","001101110111","001101111000","001101111001",
"001101111010","001101111011","001101111100","001101111101","001101111110","001101111111","001110000000","001110000001","001110000010","001110000011",
"001110000100","001110000101","001110000110","001110000111","001110001000","001110001001","001110001010","001110001011","001110001100","001110001101",
"001110001101","001110001110","001110001111","001110010000","001110010001","001110010010","001110010011","001110010100","001110010101","001110010110",
"001110010111","001110011000","001110011001","001110011010","001110011011","001110011100","001110011101","001110011110","001110011111","001110100000",
"001110100001","001110100010","001110100011","001110100100","001110100101","001110100110","001110100111","001110100111","001110101000","001110101001",
"001110101010","001110101011","001110101100","001110101101","001110101110","001110101111","001110110000","001110110001","001110110010","001110110011",
"001110110100","001110110101","001110110110","001110110111","001110111000","001110111001","001110111010","001110111011","001110111100","001110111101",
"001110111110","001110111111","001111000000","001111000001","001111000010","001111000011","001111000100","001111000100","001111000101","001111000110",
"001111000111","001111001000","001111001001","001111001010","001111001011","001111001100","001111001101","001111001110","001111001111","001111010000",
"001111010001","001111010010","001111010011","001111010100","001111010101","001111010110","001111010111","001111011000","001111011001","001111011010",
"001111011011","001111011100","001111011101","001111011110","001111011111","001111100000","001111100001","001111100010","001111100010","001111100011",
"001111100100","001111100101","001111100110","001111100111","001111101000","001111101001","001111101010","001111101011","001111101100","001111101101",
"001111101110","001111101111","001111110000","001111110001","001111110010","001111110011","001111110100","001111110101","001111110110","001111110111",
"001111111000","001111111001","001111111010","001111111011","001111111100","001111111101","001111111110","001111111111","010000000000","010000000000",
"010000000001","010000000010","010000000011","010000000100","010000000101","010000000110","010000000111","010000001000","010000001001","010000001010",
"010000001011","010000001100","010000001101","010000001110","010000001111","010000010000","010000010001","010000010010","010000010011","010000010100",
"010000010101","010000010110","010000010111","010000011000","010000011001","010000011010","010000011011","010000011100","010000011100","010000011101",
"010000011110","010000011111","010000100000","010000100001","010000100010","010000100011","010000100100","010000100101","010000100110","010000100111",
"010000101000","010000101001","010000101010","010000101011","010000101100","010000101101","010000101110","010000101111","010000110000","010000110001",
"010000110010","010000110011","010000110100","010000110101","010000110101","010000110110","010000110111","010000111000","010000111001","010000111010",
"010000111011","010000111100","010000111101","010000111110","010000111111","010001000000","010001000001","010001000010","010001000011","010001000100",
"010001000101","010001000110","010001000111","010001001000","010001001001","010001001010","010001001011","010001001100","010001001100","010001001101",
"010001001110","010001001111","010001010000","010001010001","010001010010","010001010011","010001010100","010001010101","010001010110","010001010111",
"010001011000","010001011001","010001011010","010001011011","010001011100","010001011101","010001011110","010001011111","010001100000","010001100000",
"010001100001","010001100010","010001100011","010001100100","010001100101","010001100110","010001100111","010001101000","010001101001","010001101010",
"010001101011","010001101100","010001101101","010001101110","010001101111","010001110000","010001110001","010001110010","010001110011","010001110011",
"010001110100","010001110101","010001110110","010001110111","010001111000","010001111001","010001111010","010001111011","010001111100","010001111101",
"010001111110","010001111111","010010000000","010010000001","010010000010","010010000011","010010000011","010010000100","010010000101","010010000110",
"010010000111","010010001000","010010001001","010010001010","010010001011","010010001100","010010001101","010010001110","010010001111","010010010000",
"010010010001","010010010010","010010010010","010010010011","010010010100","010010010101","010010010110","010010010111","010010011000","010010011001",
"010010011010","010010011011","010010011100","010010011101","010010011110","010010011111","010010011111","010010100000","010010100001","010010100010",
"010010100011","010010100100","010010100101","010010100110","010010100111","010010101000","010010101001","010010101010","010010101011","010010101100",
"010010101100","010010101101","010010101110","010010101111","010010110000","010010110001","010010110010","010010110011","010010110100","010010110101",
"010010110110","010010110111","010010110111","010010111000","010010111001","010010111010","010010111011","010010111100","010010111101","010010111110",
"010010111111","010011000000","010011000001","010011000010","010011000010","010011000011","010011000100","010011000101","010011000110","010011000111",
"010011001000","010011001001","010011001010","010011001011","010011001100","010011001100","010011001101","010011001110","010011001111","010011010000",
"010011010001","010011010010","010011010011","010011010100","010011010101","010011010101","010011010110","010011010111","010011011000","010011011001",
"010011011010","010011011011","010011011100","010011011101","010011011110","010011011110","010011011111","010011100000","010011100001","010011100010",
"010011100011","010011100100","010011100101","010011100110","010011100110","010011100111","010011101000","010011101001","010011101010","010011101011",
"010011101100","010011101101","010011101110","010011101110","010011101111","010011110000","010011110001","010011110010","010011110011","010011110100",
"010011110101","010011110110","010011110110","010011110111","010011111000","010011111001","010011111010","010011111011","010011111100","010011111101",
"010011111101","010011111110","010011111111","010100000000","010100000001","010100000010","010100000011","010100000100","010100000100","010100000101",
"010100000110","010100000111","010100001000","010100001001","010100001010","010100001010","010100001011","010100001100","010100001101","010100001110",
"010100001111","010100010000","010100010001","010100010001","010100010010","010100010011","010100010100","010100010101","010100010110","010100010111",
"010100010111","010100011000","010100011001","010100011010","010100011011","010100011100","010100011101","010100011101","010100011110","010100011111",
"010100100000","010100100001","010100100010","010100100010","010100100011","010100100100","010100100101","010100100110","010100100111","010100101000",
"010100101000","010100101001","010100101010","010100101011","010100101100","010100101101","010100101101","010100101110","010100101111","010100110000",
"010100110001","010100110010","010100110010","010100110011","010100110100","010100110101","010100110110","010100110111","010100110111","010100111000",
"010100111001","010100111010","010100111011","010100111100","010100111100","010100111101","010100111110","010100111111","010101000000","010101000000",
"010101000001","010101000010","010101000011","010101000100","010101000101","010101000101","010101000110","010101000111","010101001000","010101001001",
"010101001001","010101001010","010101001011","010101001100","010101001101","010101001101","010101001110","010101001111","010101010000","010101010001",
"010101010010","010101010010","010101010011","010101010100","010101010101","010101010110","010101010110","010101010111","010101011000","010101011001",
"010101011001","010101011010","010101011011","010101011100","010101011101","010101011101","010101011110","010101011111","010101100000","010101100001",
"010101100001","010101100010","010101100011","010101100100","010101100101","010101100101","010101100110","010101100111","010101101000","010101101000",
"010101101001","010101101010","010101101011","010101101100","010101101100","010101101101","010101101110","010101101111","010101101111","010101110000",
"010101110001","010101110010","010101110010","010101110011","010101110100","010101110101","010101110110","010101110110","010101110111","010101111000",
"010101111001","010101111001","010101111010","010101111011","010101111100","010101111100","010101111101","010101111110","010101111111","010101111111",
"010110000000","010110000001","010110000010","010110000010","010110000011","010110000100","010110000101","010110000101","010110000110","010110000111",
"010110001000","010110001000","010110001001","010110001010","010110001011","010110001011","010110001100","010110001101","010110001101","010110001110",
"010110001111","010110010000","010110010000","010110010001","010110010010","010110010011","010110010011","010110010100","010110010101","010110010101",
"010110010110","010110010111","010110011000","010110011000","010110011001","010110011010","010110011010","010110011011","010110011100","010110011101",
"010110011101","010110011110","010110011111","010110011111","010110100000","010110100001","010110100010","010110100010","010110100011","010110100100",
"010110100100","010110100101","010110100110","010110100110","010110100111","010110101000","010110101001","010110101001","010110101010","010110101011",
"010110101011","010110101100","010110101101","010110101101","010110101110","010110101111","010110101111","010110110000","010110110001","010110110001",
"010110110010","010110110011","010110110100","010110110100","010110110101","010110110110","010110110110","010110110111","010110111000","010110111000",
"010110111001","010110111010","010110111010","010110111011","010110111100","010110111100","010110111101","010110111110","010110111110","010110111111",
"010111000000","010111000000","010111000001","010111000001","010111000010","010111000011","010111000011","010111000100","010111000101","010111000101",
"010111000110","010111000111","010111000111","010111001000","010111001001","010111001001","010111001010","010111001011","010111001011","010111001100",
"010111001100","010111001101","010111001110","010111001110","010111001111","010111010000","010111010000","010111010001","010111010001","010111010010",
"010111010011","010111010011","010111010100","010111010101","010111010101","010111010110","010111010110","010111010111","010111011000","010111011000",
"010111011001","010111011010","010111011010","010111011011","010111011011","010111011100","010111011101","010111011101","010111011110","010111011110",
"010111011111","010111100000","010111100000","010111100001","010111100001","010111100010","010111100011","010111100011","010111100100","010111100100",
"010111100101","010111100101","010111100110","010111100111","010111100111","010111101000","010111101000","010111101001","010111101010","010111101010",
"010111101011","010111101011","010111101100","010111101100","010111101101","010111101110","010111101110","010111101111","010111101111","010111110000",
"010111110000","010111110001","010111110010","010111110010","010111110011","010111110011","010111110100","010111110100","010111110101","010111110101",
"010111110110","010111110110","010111110111","010111111000","010111111000","010111111001","010111111001","010111111010","010111111010","010111111011",
"010111111011","010111111100","010111111100","010111111101","010111111110","010111111110","010111111111","010111111111","011000000000","011000000000",
"011000000001","011000000001","011000000010","011000000010","011000000011","011000000011","011000000100","011000000100","011000000101","011000000101",
"011000000110","011000000110","011000000111","011000000111","011000001000","011000001000","011000001001","011000001001","011000001010","011000001010",
"011000001011","011000001011","011000001100","011000001100","011000001101","011000001101","011000001110","011000001110","011000001111","011000001111",
"011000010000","011000010000","011000010001","011000010001","011000010010","011000010010","011000010011","011000010011","011000010100","011000010100",
"011000010101","011000010101","011000010110","011000010110","011000010111","011000010111","011000010111","011000011000","011000011000","011000011001",
"011000011001","011000011010","011000011010","011000011011","011000011011","011000011100","011000011100","011000011100","011000011101","011000011101",
"011000011110","011000011110","011000011111","011000011111","011000100000","011000100000","011000100000","011000100001","011000100001","011000100010",
"011000100010","011000100011","011000100011","011000100011","011000100100","011000100100","011000100101","011000100101","011000100110","011000100110",
"011000100110","011000100111","011000100111","011000101000","011000101000","011000101001","011000101001","011000101001","011000101010","011000101010",
"011000101011","011000101011","011000101011","011000101100","011000101100","011000101101","011000101101","011000101101","011000101110","011000101110",
"011000101111","011000101111","011000101111","011000110000","011000110000","011000110000","011000110001","011000110001","011000110010","011000110010",
"011000110010","011000110011","011000110011","011000110011","011000110100","011000110100","011000110101","011000110101","011000110101","011000110110",
"011000110110","011000110110","011000110111","011000110111","011000110111","011000111000","011000111000","011000111001","011000111001","011000111001",
"011000111010","011000111010","011000111010","011000111011","011000111011","011000111011","011000111100","011000111100","011000111100","011000111101",
"011000111101","011000111101","011000111110","011000111110","011000111110","011000111111","011000111111","011000111111","011001000000","011001000000",
"011001000000","011001000001","011001000001","011001000001","011001000001","011001000010","011001000010","011001000010","011001000011","011001000011",
"011001000011","011001000100","011001000100","011001000100","011001000101","011001000101","011001000101","011001000101","011001000110","011001000110",
"011001000110","011001000111","011001000111","011001000111","011001000111","011001001000","011001001000","011001001000","011001001001","011001001001",
"011001001001","011001001001","011001001010","011001001010","011001001010","011001001010","011001001011","011001001011","011001001011","011001001011",
"011001001100","011001001100","011001001100","011001001100","011001001101","011001001101","011001001101","011001001101","011001001110","011001001110",
"011001001110","011001001110","011001001111","011001001111","011001001111","011001001111","011001010000","011001010000","011001010000","011001010000",
"011001010001","011001010001","011001010001","011001010001","011001010001","011001010010","011001010010","011001010010","011001010010","011001010011",
"011001010011","011001010011","011001010011","011001010011","011001010100","011001010100","011001010100","011001010100","011001010100","011001010101",
"011001010101","011001010101","011001010101","011001010101","011001010110","011001010110","011001010110","011001010110","011001010110","011001010111",
"011001010111","011001010111","011001010111","011001010111","011001010111","011001011000","011001011000","011001011000","011001011000","011001011000",
"011001011001","011001011001","011001011001","011001011001","011001011001","011001011001","011001011001","011001011010","011001011010","011001011010",
"011001011010","011001011010","011001011010","011001011011","011001011011","011001011011","011001011011","011001011011","011001011011","011001011011",
"011001011100","011001011100","011001011100","011001011100","011001011100","011001011100","011001011100","011001011100","011001011101","011001011101",
"011001011101","011001011101","011001011101","011001011101","011001011101","011001011101","011001011110","011001011110","011001011110","011001011110",
"011001011110","011001011110","011001011110","011001011110","011001011110","011001011110","011001011111","011001011111","011001011111","011001011111",
"011001011111","011001011111","011001011111","011001011111","011001011111","011001011111","011001011111","011001100000","011001100000","011001100000",
"011001100000","011001100000","011001100000","011001100000","011001100000","011001100000","011001100000","011001100000","011001100000","011001100000",
"011001100000","011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100001",
"011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100001",
"011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100010",
"011001100010","011001100010","011001100010","011001100010","011001100010","011001100010","011001100010","011001100010","011001100010","011001100010",
"011001100010","011001100010","011001100010","011001100010","011001100010","011001100010","011001100010","011001100010","011001100001","011001100001",
"011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100001",
"011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100001",
"011001100001","011001100001","011001100001","011001100001","011001100001","011001100001","011001100000","011001100000","011001100000","011001100000",
"011001100000","011001100000","011001100000","011001100000","011001100000","011001100000","011001100000","011001100000","011001100000","011001100000",
"011001011111","011001011111","011001011111","011001011111","011001011111","011001011111","011001011111","011001011111","011001011111","011001011111",
"011001011111","011001011110","011001011110","011001011110","011001011110","011001011110","011001011110","011001011110","011001011110","011001011110",
"011001011110","011001011101","011001011101","011001011101","011001011101","011001011101","011001011101","011001011101","011001011101","011001011100",
"011001011100","011001011100","011001011100","011001011100","011001011100","011001011100","011001011100","011001011011","011001011011","011001011011",
"011001011011","011001011011","011001011011","011001011011","011001011010","011001011010","011001011010","011001011010","011001011010","011001011010",
"011001011001","011001011001","011001011001","011001011001","011001011001","011001011001","011001011001","011001011000","011001011000","011001011000",
"011001011000","011001011000","011001010111","011001010111","011001010111","011001010111","011001010111","011001010111","011001010110","011001010110",
"011001010110","011001010110","011001010110","011001010101","011001010101","011001010101","011001010101","011001010101","011001010100","011001010100",
"011001010100","011001010100","011001010100","011001010011","011001010011","011001010011","011001010011","011001010011","011001010010","011001010010",
"011001010010","011001010010","011001010001","011001010001","011001010001","011001010001","011001010001","011001010000","011001010000","011001010000",
"011001010000","011001001111","011001001111","011001001111","011001001111","011001001110","011001001110","011001001110","011001001110","011001001101",
"011001001101","011001001101","011001001101","011001001100","011001001100","011001001100","011001001100","011001001011","011001001011","011001001011",
"011001001011","011001001010","011001001010","011001001010","011001001010","011001001001","011001001001","011001001001","011001001001","011001001000",
"011001001000","011001001000","011001000111","011001000111","011001000111","011001000111","011001000110","011001000110","011001000110","011001000101",
"011001000101","011001000101","011001000101","011001000100","011001000100","011001000100","011001000011","011001000011","011001000011","011001000010",
"011001000010","011001000010","011001000001","011001000001","011001000001","011001000001","011001000000","011001000000","011001000000","011000111111",
"011000111111","011000111111","011000111110","011000111110","011000111110","011000111101","011000111101","011000111101","011000111100","011000111100",
"011000111100","011000111011","011000111011","011000111011","011000111010","011000111010","011000111010","011000111001","011000111001","011000111001",
"011000111000","011000111000","011000110111","011000110111","011000110111","011000110110","011000110110","011000110110","011000110101","011000110101",
"011000110101","011000110100","011000110100","011000110011","011000110011","011000110011","011000110010","011000110010","011000110010","011000110001",
"011000110001","011000110000","011000110000","011000110000","011000101111","011000101111","011000101111","011000101110","011000101110","011000101101",
"011000101101","011000101101","011000101100","011000101100","011000101011","011000101011","011000101011","011000101010","011000101010","011000101001",
"011000101001","011000101001","011000101000","011000101000","011000100111","011000100111","011000100110","011000100110","011000100110","011000100101",
"011000100101","011000100100","011000100100","011000100011","011000100011","011000100011","011000100010","011000100010","011000100001","011000100001",
"011000100000","011000100000","011000100000","011000011111","011000011111","011000011110","011000011110","011000011101","011000011101","011000011100",
"011000011100","011000011100","011000011011","011000011011","011000011010","011000011010","011000011001","011000011001","011000011000","011000011000",
"011000010111","011000010111","011000010111","011000010110","011000010110","011000010101","011000010101","011000010100","011000010100","011000010011",
"011000010011","011000010010","011000010010","011000010001","011000010001","011000010000","011000010000","011000001111","011000001111","011000001110",
"011000001110","011000001101","011000001101","011000001100","011000001100","011000001011","011000001011","011000001010","011000001010","011000001001",
"011000001001","011000001000","011000001000","011000000111","011000000111","011000000110","011000000110","011000000101","011000000101","011000000100",
"011000000100","011000000011","011000000011","011000000010","011000000010","011000000001","011000000001","011000000000","011000000000","010111111111",
"010111111111","010111111110","010111111110","010111111101","010111111100","010111111100","010111111011","010111111011","010111111010","010111111010",
"010111111001","010111111001","010111111000","010111111000","010111110111","010111110110","010111110110","010111110101","010111110101","010111110100",
"010111110100","010111110011","010111110011","010111110010","010111110010","010111110001","010111110000","010111110000","010111101111","010111101111",
"010111101110","010111101110","010111101101","010111101100","010111101100","010111101011","010111101011","010111101010","010111101010","010111101001",
"010111101000","010111101000","010111100111","010111100111","010111100110","010111100101","010111100101","010111100100","010111100100","010111100011",
"010111100011","010111100010","010111100001","010111100001","010111100000","010111100000","010111011111","010111011110","010111011110","010111011101",
"010111011101","010111011100","010111011011","010111011011","010111011010","010111011010","010111011001","010111011000","010111011000","010111010111",
"010111010110","010111010110","010111010101","010111010101","010111010100","010111010011","010111010011","010111010010","010111010001","010111010001",
"010111010000","010111010000","010111001111","010111001110","010111001110","010111001101","010111001100","010111001100","010111001011","010111001011",
"010111001010","010111001001","010111001001","010111001000","010111000111","010111000111","010111000110","010111000101","010111000101","010111000100",
"010111000011","010111000011","010111000010","010111000001","010111000001","010111000000","010111000000","010110111111","010110111110","010110111110",
"010110111101","010110111100","010110111100","010110111011","010110111010","010110111010","010110111001","010110111000","010110111000","010110110111",
"010110110110","010110110110","010110110101","010110110100","010110110100","010110110011","010110110010","010110110001","010110110001","010110110000",
"010110101111","010110101111","010110101110","010110101101","010110101101","010110101100","010110101011","010110101011","010110101010","010110101001",
"010110101001","010110101000","010110100111","010110100110","010110100110","010110100101","010110100100","010110100100","010110100011","010110100010",
"010110100010","010110100001","010110100000","010110011111","010110011111","010110011110","010110011101","010110011101","010110011100","010110011011",
"010110011010","010110011010","010110011001","010110011000","010110011000","010110010111","010110010110","010110010101","010110010101","010110010100",
"010110010011","010110010011","010110010010","010110010001","010110010000","010110010000","010110001111","010110001110","010110001101","010110001101",
"010110001100","010110001011","010110001011","010110001010","010110001001","010110001000","010110001000","010110000111","010110000110","010110000101",
"010110000101","010110000100","010110000011","010110000010","010110000010","010110000001","010110000000","010101111111","010101111111","010101111110",
"010101111101","010101111100","010101111100","010101111011","010101111010","010101111001","010101111001","010101111000","010101110111","010101110110",
"010101110110","010101110101","010101110100","010101110011","010101110010","010101110010","010101110001","010101110000","010101101111","010101101111",
"010101101110","010101101101","010101101100","010101101100","010101101011","010101101010","010101101001","010101101000","010101101000","010101100111",
"010101100110","010101100101","010101100101","010101100100","010101100011","010101100010","010101100001","010101100001","010101100000","010101011111",
"010101011110","010101011101","010101011101","010101011100","010101011011","010101011010","010101011001","010101011001","010101011000","010101010111",
"010101010110","010101010110","010101010101","010101010100","010101010011","010101010010","010101010010","010101010001","010101010000","010101001111",
"010101001110","010101001101","010101001101","010101001100","010101001011","010101001010","010101001001","010101001001","010101001000","010101000111",
"010101000110","010101000101","010101000101","010101000100","010101000011","010101000010","010101000001","010101000000","010101000000","010100111111",
"010100111110","010100111101","010100111100","010100111100","010100111011","010100111010","010100111001","010100111000","010100110111","010100110111",
"010100110110","010100110101","010100110100","010100110011","010100110010","010100110010","010100110001","010100110000","010100101111","010100101110",
"010100101101","010100101101","010100101100","010100101011","010100101010","010100101001","010100101000","010100101000","010100100111","010100100110",
"010100100101","010100100100","010100100011","010100100010","010100100010","010100100001","010100100000","010100011111","010100011110","010100011101",
"010100011101","010100011100","010100011011","010100011010","010100011001","010100011000","010100010111","010100010111","010100010110","010100010101",
"010100010100","010100010011","010100010010","010100010001","010100010001","010100010000","010100001111","010100001110","010100001101","010100001100",
"010100001011","010100001010","010100001010","010100001001","010100001000","010100000111","010100000110","010100000101","010100000100","010100000100",
"010100000011","010100000010","010100000001","010100000000","010011111111","010011111110","010011111101","010011111101","010011111100","010011111011",
"010011111010","010011111001","010011111000","010011110111","010011110110","010011110110","010011110101","010011110100","010011110011","010011110010",
"010011110001","010011110000","010011101111","010011101110","010011101110","010011101101","010011101100","010011101011","010011101010","010011101001",
"010011101000","010011100111","010011100110","010011100110","010011100101","010011100100","010011100011","010011100010","010011100001","010011100000",
"010011011111","010011011110","010011011110","010011011101","010011011100","010011011011","010011011010","010011011001","010011011000","010011010111",
"010011010110","010011010101","010011010101","010011010100","010011010011","010011010010","010011010001","010011010000","010011001111","010011001110",
"010011001101","010011001100","010011001100","010011001011","010011001010","010011001001","010011001000","010011000111","010011000110","010011000101",
"010011000100","010011000011","010011000010","010011000010","010011000001","010011000000","010010111111","010010111110","010010111101","010010111100",
"010010111011","010010111010","010010111001","010010111000","010010110111","010010110111","010010110110","010010110101","010010110100","010010110011",
"010010110010","010010110001","010010110000","010010101111","010010101110","010010101101","010010101100","010010101100","010010101011","010010101010",
"010010101001","010010101000","010010100111","010010100110","010010100101","010010100100","010010100011","010010100010","010010100001","010010100000",
"010010011111","010010011111","010010011110","010010011101","010010011100","010010011011","010010011010","010010011001","010010011000","010010010111",
"010010010110","010010010101","010010010100","010010010011","010010010010","010010010010","010010010001","010010010000","010010001111","010010001110",
"010010001101","010010001100","010010001011","010010001010","010010001001","010010001000","010010000111","010010000110","010010000101","010010000100",
"010010000011","010010000011","010010000010","010010000001","010010000000","010001111111","010001111110","010001111101","010001111100","010001111011",
"010001111010","010001111001","010001111000","010001110111","010001110110","010001110101","010001110100","010001110011","010001110011","010001110010",
"010001110001","010001110000","010001101111","010001101110","010001101101","010001101100","010001101011","010001101010","010001101001","010001101000",
"010001100111","010001100110","010001100101","010001100100","010001100011","010001100010","010001100001","010001100000","010001100000","010001011111",
"010001011110","010001011101","010001011100","010001011011","010001011010","010001011001","010001011000","010001010111","010001010110","010001010101",
"010001010100","010001010011","010001010010","010001010001","010001010000","010001001111","010001001110","010001001101","010001001100","010001001100",
"010001001011","010001001010","010001001001","010001001000","010001000111","010001000110","010001000101","010001000100","010001000011","010001000010",
"010001000001","010001000000","010000111111","010000111110","010000111101","010000111100","010000111011","010000111010","010000111001","010000111000",
"010000110111","010000110110","010000110101","010000110101","010000110100","010000110011","010000110010","010000110001","010000110000","010000101111",
"010000101110","010000101101","010000101100","010000101011","010000101010","010000101001","010000101000","010000100111","010000100110","010000100101",
"010000100100","010000100011","010000100010","010000100001","010000100000","010000011111","010000011110","010000011101","010000011100","010000011100",
"010000011011","010000011010","010000011001","010000011000","010000010111","010000010110","010000010101","010000010100","010000010011","010000010010",
"010000010001","010000010000","010000001111","010000001110","010000001101","010000001100","010000001011","010000001010","010000001001","010000001000",
"010000000111","010000000110","010000000101","010000000100","010000000011","010000000010","010000000001","010000000000","010000000000","001111111111",
"001111111110","001111111101","001111111100","001111111011","001111111010","001111111001","001111111000","001111110111","001111110110","001111110101",
"001111110100","001111110011","001111110010","001111110001","001111110000","001111101111","001111101110","001111101101","001111101100","001111101011",
"001111101010","001111101001","001111101000","001111100111","001111100110","001111100101","001111100100","001111100011","001111100010","001111100010",
"001111100001","001111100000","001111011111","001111011110","001111011101","001111011100","001111011011","001111011010","001111011001","001111011000",
"001111010111","001111010110","001111010101","001111010100","001111010011","001111010010","001111010001","001111010000","001111001111","001111001110",
"001111001101","001111001100","001111001011","001111001010","001111001001","001111001000","001111000111","001111000110","001111000101","001111000100",
"001111000100","001111000011","001111000010","001111000001","001111000000","001110111111","001110111110","001110111101","001110111100","001110111011",
"001110111010","001110111001","001110111000","001110110111","001110110110","001110110101","001110110100","001110110011","001110110010","001110110001",
"001110110000","001110101111","001110101110","001110101101","001110101100","001110101011","001110101010","001110101001","001110101000","001110100111",
"001110100111","001110100110","001110100101","001110100100","001110100011","001110100010","001110100001","001110100000","001110011111","001110011110",
"001110011101","001110011100","001110011011","001110011010","001110011001","001110011000","001110010111","001110010110","001110010101","001110010100",
"001110010011","001110010010","001110010001","001110010000","001110001111","001110001110","001110001101","001110001101","001110001100","001110001011",
"001110001010","001110001001","001110001000","001110000111","001110000110","001110000101","001110000100","001110000011","001110000010","001110000001",
"001110000000","001101111111","001101111110","001101111101","001101111100","001101111011","001101111010","001101111001","001101111000","001101110111",
"001101110110","001101110110","001101110101","001101110100","001101110011","001101110010","001101110001","001101110000","001101101111","001101101110",
"001101101101","001101101100","001101101011","001101101010","001101101001","001101101000","001101100111","001101100110","001101100101","001101100100",
"001101100011","001101100010","001101100001","001101100000","001101100000","001101011111","001101011110","001101011101","001101011100","001101011011",
"001101011010","001101011001","001101011000","001101010111","001101010110","001101010101","001101010100","001101010011","001101010010","001101010001",
"001101010000","001101001111","001101001110","001101001101","001101001101","001101001100","001101001011","001101001010","001101001001","001101001000",
"001101000111","001101000110","001101000101","001101000100","001101000011","001101000010","001101000001","001101000000","001100111111","001100111110",
"001100111101","001100111100","001100111100","001100111011","001100111010","001100111001","001100111000","001100110111","001100110110","001100110101",
"001100110100","001100110011","001100110010","001100110001","001100110000","001100101111","001100101110","001100101101","001100101100","001100101100",
"001100101011","001100101010","001100101001","001100101000","001100100111","001100100110","001100100101","001100100100","001100100011","001100100010",
"001100100001","001100100000","001100011111","001100011110","001100011101","001100011101","001100011100","001100011011","001100011010","001100011001",
"001100011000","001100010111","001100010110","001100010101","001100010100","001100010011","001100010010","001100010001","001100010000","001100010000",
"001100001111","001100001110","001100001101","001100001100","001100001011","001100001010","001100001001","001100001000","001100000111","001100000110",
"001100000101","001100000100","001100000100","001100000011","001100000010","001100000001","001100000000","001011111111","001011111110","001011111101",
"001011111100","001011111011","001011111010","001011111001","001011111000","001011111000","001011110111","001011110110","001011110101","001011110100",
"001011110011","001011110010","001011110001","001011110000","001011101111","001011101110","001011101101","001011101101","001011101100","001011101011",
"001011101010","001011101001","001011101000","001011100111","001011100110","001011100101","001011100100","001011100011","001011100011","001011100010",
"001011100001","001011100000","001011011111","001011011110","001011011101","001011011100","001011011011","001011011010","001011011001","001011011001",
"001011011000","001011010111","001011010110","001011010101","001011010100","001011010011","001011010010","001011010001","001011010000","001011010000",
"001011001111","001011001110","001011001101","001011001100","001011001011","001011001010","001011001001","001011001000","001011000111","001011000111",
"001011000110","001011000101","001011000100","001011000011","001011000010","001011000001","001011000000","001010111111","001010111110","001010111110",
"001010111101","001010111100","001010111011","001010111010","001010111001","001010111000","001010110111","001010110110","001010110110","001010110101",
"001010110100","001010110011","001010110010","001010110001","001010110000","001010101111","001010101111","001010101110","001010101101","001010101100",
"001010101011","001010101010","001010101001","001010101000","001010100111","001010100111","001010100110","001010100101","001010100100","001010100011",
"001010100010","001010100001","001010100000","001010100000","001010011111","001010011110","001010011101","001010011100","001010011011","001010011010",
"001010011001","001010011001","001010011000","001010010111","001010010110","001010010101","001010010100","001010010011","001010010011","001010010010",
"001010010001","001010010000","001010001111","001010001110","001010001101","001010001100","001010001100","001010001011","001010001010","001010001001",
"001010001000","001010000111","001010000110","001010000110","001010000101","001010000100","001010000011","001010000010","001010000001","001010000000",
"001010000000","001001111111","001001111110","001001111101","001001111100","001001111011","001001111010","001001111010","001001111001","001001111000",
"001001110111","001001110110","001001110101","001001110100","001001110100","001001110011","001001110010","001001110001","001001110000","001001101111",
"001001101111","001001101110","001001101101","001001101100","001001101011","001001101010","001001101001","001001101001","001001101000","001001100111",
"001001100110","001001100101","001001100100","001001100100","001001100011","001001100010","001001100001","001001100000","001001011111","001001011111",
"001001011110","001001011101","001001011100","001001011011","001001011010","001001011010","001001011001","001001011000","001001010111","001001010110",
"001001010101","001001010101","001001010100","001001010011","001001010010","001001010001","001001010000","001001010000","001001001111","001001001110",
"001001001101","001001001100","001001001100","001001001011","001001001010","001001001001","001001001000","001001000111","001001000111","001001000110",
"001001000101","001001000100","001001000011","001001000011","001001000010","001001000001","001001000000","001000111111","001000111110","001000111110",
"001000111101","001000111100","001000111011","001000111010","001000111010","001000111001","001000111000","001000110111","001000110110","001000110110",
"001000110101","001000110100","001000110011","001000110010","001000110010","001000110001","001000110000","001000101111","001000101110","001000101110",
"001000101101","001000101100","001000101011","001000101010","001000101010","001000101001","001000101000","001000100111","001000100110","001000100110",
"001000100101","001000100100","001000100011","001000100010","001000100010","001000100001","001000100000","001000011111","001000011111","001000011110",
"001000011101","001000011100","001000011011","001000011011","001000011010","001000011001","001000011000","001000010111","001000010111","001000010110",
"001000010101","001000010100","001000010100","001000010011","001000010010","001000010001","001000010000","001000010000","001000001111","001000001110",
"001000001101","001000001101","001000001100","001000001011","001000001010","001000001001","001000001001","001000001000","001000000111","001000000110",
"001000000110","001000000101","001000000100","001000000011","001000000011","001000000010","001000000001","001000000000","001000000000","000111111111",
"000111111110","000111111101","000111111100","000111111100","000111111011","000111111010","000111111001","000111111001","000111111000","000111110111",
"000111110110","000111110110","000111110101","000111110100","000111110011","000111110011","000111110010","000111110001","000111110000","000111110000",
"000111101111","000111101110","000111101101","000111101101","000111101100","000111101011","000111101010","000111101010","000111101001","000111101000",
"000111100111","000111100111","000111100110","000111100101","000111100101","000111100100","000111100011","000111100010","000111100010","000111100001",
"000111100000","000111011111","000111011111","000111011110","000111011101","000111011100","000111011100","000111011011","000111011010","000111011010",
"000111011001","000111011000","000111010111","000111010111","000111010110","000111010101","000111010100","000111010100","000111010011","000111010010",
"000111010010","000111010001","000111010000","000111001111","000111001111","000111001110","000111001101","000111001101","000111001100","000111001011",
"000111001010","000111001010","000111001001","000111001000","000111001000","000111000111","000111000110","000111000101","000111000101","000111000100",
"000111000011","000111000011","000111000010","000111000001","000111000000","000111000000","000110111111","000110111110","000110111110","000110111101",
"000110111100","000110111100","000110111011","000110111010","000110111001","000110111001","000110111000","000110110111","000110110111","000110110110",
"000110110101","000110110101","000110110100","000110110011","000110110010","000110110010","000110110001","000110110000","000110110000","000110101111",
"000110101110","000110101110","000110101101","000110101100","000110101100","000110101011","000110101010","000110101010","000110101001","000110101000",
"000110101000","000110100111","000110100110","000110100101","000110100101","000110100100","000110100011","000110100011","000110100010","000110100001",
"000110100001","000110100000","000110011111","000110011111","000110011110","000110011101","000110011101","000110011100","000110011011","000110011011",
"000110011010","000110011001","000110011001","000110011000","000110010111","000110010111","000110010110","000110010101","000110010101","000110010100",
"000110010011","000110010011","000110010010","000110010001","000110010001","000110010000","000110001111","000110001111","000110001110","000110001110",
"000110001101","000110001100","000110001100","000110001011","000110001010","000110001010","000110001001","000110001000","000110001000","000110000111",
"000110000110","000110000110","000110000101","000110000100","000110000100","000110000011","000110000011","000110000010","000110000001","000110000001",
"000110000000","000101111111","000101111111","000101111110","000101111101","000101111101","000101111100","000101111100","000101111011","000101111010",
"000101111010","000101111001","000101111000","000101111000","000101110111","000101110110","000101110110","000101110101","000101110101","000101110100",
"000101110011","000101110011","000101110010","000101110001","000101110001","000101110000","000101110000","000101101111","000101101110","000101101110",
"000101101101","000101101100","000101101100","000101101011","000101101011","000101101010","000101101001","000101101001","000101101000","000101101000",
"000101100111","000101100110","000101100110","000101100101","000101100101","000101100100","000101100011","000101100011","000101100010","000101100001",
"000101100001","000101100000","000101100000","000101011111","000101011110","000101011110","000101011101","000101011101","000101011100","000101011011",
"000101011011","000101011010","000101011010","000101011001","000101011001","000101011000","000101010111","000101010111","000101010110","000101010110",
"000101010101","000101010100","000101010100","000101010011","000101010011","000101010010","000101010001","000101010001","000101010000","000101010000",
"000101001111","000101001111","000101001110","000101001101","000101001101","000101001100","000101001100","000101001011","000101001010","000101001010",
"000101001001","000101001001","000101001000","000101001000","000101000111","000101000110","000101000110","000101000101","000101000101","000101000100",
"000101000100","000101000011","000101000010","000101000010","000101000001","000101000001","000101000000","000101000000","000100111111","000100111110",
"000100111110","000100111101","000100111101","000100111100","000100111100","000100111011","000100111011","000100111010","000100111001","000100111001",
"000100111000","000100111000","000100110111","000100110111","000100110110","000100110110","000100110101","000100110100","000100110100","000100110011",
"000100110011","000100110010","000100110010","000100110001","000100110001","000100110000","000100110000","000100101111","000100101110","000100101110",
"000100101101","000100101101","000100101100","000100101100","000100101011","000100101011","000100101010","000100101010","000100101001","000100101000",
"000100101000","000100100111","000100100111","000100100110","000100100110","000100100101","000100100101","000100100100","000100100100","000100100011",
"000100100011","000100100010","000100100010","000100100001","000100100001","000100100000","000100011111","000100011111","000100011110","000100011110",
"000100011101","000100011101","000100011100","000100011100","000100011011","000100011011","000100011010","000100011010","000100011001","000100011001",
"000100011000","000100011000","000100010111","000100010111","000100010110","000100010110","000100010101","000100010101","000100010100","000100010100",
"000100010011","000100010011","000100010010","000100010010","000100010001","000100010001","000100010000","000100010000","000100001111","000100001111",
"000100001110","000100001110","000100001101","000100001101","000100001100","000100001100","000100001011","000100001011","000100001010","000100001010",
"000100001001","000100001001","000100001000","000100001000","000100000111","000100000111","000100000110","000100000110","000100000101","000100000101",
"000100000100","000100000100","000100000011","000100000011","000100000010","000100000010","000100000001","000100000001","000100000000","000100000000",
"000011111111","000011111111","000011111110","000011111110","000011111101","000011111101","000011111100","000011111100","000011111100","000011111011",
"000011111011","000011111010","000011111010","000011111001","000011111001","000011111000","000011111000","000011110111","000011110111","000011110110",
"000011110110","000011110101","000011110101","000011110100","000011110100","000011110100","000011110011","000011110011","000011110010","000011110010",
"000011110001","000011110001","000011110000","000011110000","000011101111","000011101111","000011101110","000011101110","000011101110","000011101101",
"000011101101","000011101100","000011101100","000011101011","000011101011","000011101010","000011101010","000011101001","000011101001","000011101001",
"000011101000","000011101000","000011100111","000011100111","000011100110","000011100110","000011100101","000011100101","000011100101","000011100100",
"000011100100","000011100011","000011100011","000011100010","000011100010","000011100001","000011100001","000011100001","000011100000","000011100000",
"000011011111","000011011111","000011011110","000011011110","000011011110","000011011101");
	begin  
		process(address)
		begin
			window_val <= window_lut(to_integer(unsigned(address)));	
		end process;
end behavioral;