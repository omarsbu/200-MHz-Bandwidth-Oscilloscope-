library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_17_strings_slv is
  generic (
    STR_LEN   : natural := 16;   -- all strings are 16 chars
    STR_COUNT : natural := 17    -- total strings
  );
  port (
    clk    : in  std_logic;
    addr   : in  std_logic_vector(8 downto 0);  -- 0..271 (9 bits)
    o_char : out std_logic_vector(6 downto 0)   -- 7-bit ASCII
  );
end entity;

architecture rtl of rom_17_strings_slv is

  constant ROM_SIZE : natural := STR_LEN * STR_COUNT;

  -- Flattened ROM as character array
  type rom_type is array(0 to ROM_SIZE-1) of character;

  constant CHAR_ROM : rom_type := (
    -- str1: "100mV/DIV       "
     0=>'1',1=>'0',2=>'0',3=>'m',4=>'V',5=>'/',6=>'D',7=>'I',
     8=>'V',9=>' ',10=>' ',11=>' ',12=>' ',13=>' ',14=>' ',15=>' ',
    -- str2: "100us/DIV       "
    16=>'1',17=>'0',18=>'0',19=>'u',20=>'s',21=>'/',22=>'D',23=>'I',
    24=>'V',25=>' ',26=>' ',27=>' ',28=>' ',29=>' ',30=>' ',31=>' ',
    -- str3: "Delay: 100us    "
    32=>'D',33=>'e',34=>'l',35=>'a',36=>'y',37=>':',38=>' ',39=>'1',
    40=>'0',41=>'0',42=>'u',43=>'s',44=>' ',45=>' ',46=>' ',47=>' ',
    -- str4: "TRG LVL: 100mV  "
    48=>'T',49=>'R',50=>'G',51=>' ',52=>'L',53=>'V',54=>'L',55=>':',
    56=>' ',57=>'1',58=>'0',59=>'0',60=>'m',61=>'V',62=>' ',63=>' ',
    -- str5: "(RISING)        "
    64=>'(',65=>'R',66=>'I',67=>'S',68=>'I',69=>'N',70=>'G',71=>')',
    72=>' ',73=>' ',74=>' ',75=>' ',76=>' ',77=>' ',78=>' ',79=>' ',
    -- str6: "100MSa/s        "
    80=>'1',81=>'0',82=>'0',83=>'M',84=>'S',85=>'a',86=>'/',87=>'s',
    88=>' ',89=>' ',90=>' ',91=>' ',92=>' ',93=>' ',94=>' ',95=>' ',
    -- str7: "Freq: 100MHz    "
    96=>'F',97=>'r',98=>'e',99=>'q',100=>':',101=>' ',102=>'1',103=>'0',
   104=>'0',105=>'M',106=>'H',107=>'z',108=>' ',109=>' ',110=>' ',111=>' ',
    -- str8: "V(max): 100mV   "
   112=>'V',113=>'(',114=>'m',115=>'a',116=>'x',117=>')',118=>':',
   119=>' ',120=>'1',121=>'0',122=>'0',123=>'m',124=>'V',125=>' ',126=>' ',127=>' ',
    -- str9: "V(min): 100mV   "
   128=>'V',129=>'(',130=>'m',131=>'i',132=>'n',133=>')',134=>':',
   135=>' ',136=>'1',137=>'0',138=>'0',139=>'m',140=>'V',141=>' ',142=>' ',143=>' ',
    -- str10: "V(avg): 100mV   "
   144=>'V',145=>'(',146=>'a',147=>'v',148=>'g',149=>')',150=>':',
   151=>' ',152=>'1',153=>'0',154=>'0',155=>'m',156=>'V',157=>' ',158=>' ',159=>' ',
    -- str11: "V(p-p): 100mV   "
   160=>'V',161=>'(',162=>'p',163=>'-',164=>'p',165=>')',166=>':',
   167=>' ',168=>'1',169=>'0',170=>'0',171=>'m',172=>'V',173=>' ',174=>' ',175=>' ',
    -- str12: "X1: 100us       "
   176=>'X',177=>'1',178=>':',179=>' ',180=>'1',181=>'0',182=>'0',183=>'u',
   184=>'s',185=>' ',186=>' ',187=>' ',188=>' ',189=>' ',190=>' ',191=>' ',
    -- str13: "X2: 100us       "
   192=>'X',193=>'2',194=>':',195=>' ',196=>'1',197=>'0',198=>'0',199=>'u',
   200=>'s',201=>' ',202=>' ',203=>' ',204=>' ',205=>' ',206=>' ',207=>' ',
    -- str14: "Y1: 100mV       "
   208=>'Y',209=>'1',210=>':',211=>' ',212=>'1',213=>'0',214=>'0',215=>'m',
   216=>'V',217=>' ',218=>' ',219=>' ',220=>' ',221=>' ',222=>' ',223=>' ',
    -- str15: "Y2: 100mV       "
   224=>'Y',225=>'2',226=>':',227=>' ',228=>'1',229=>'0',230=>'0',231=>'m',
   232=>'V',233=>' ',234=>' ',235=>' ',236=>' ',237=>' ',238=>' ',239=>' ',
    -- str16: "(X2-X1): 100us  "
   240=>'(',241=>'X',242=>'2',243=>'-',244=>'X',245=>'1',246=>')',247=>':',
   248=>' ',249=>'1',250=>'0',251=>'0',252=>'u',253=>'s',254=>' ',255=>' ',
    -- str17: "(Y2-Y1): 100mV  "
   256=>'(',257=>'Y',258=>'2',259=>'-',260=>'Y',261=>'1',262=>')',263=>':',
   264=>' ',265=>'1',266=>'0',267=>'0',268=>'m',269=>'V',270=>' ',271=>' '
  );

  -- Convert character to 7-bit SLV
  function char_to_slv(c: character) return std_logic_vector is
  begin
    return std_logic_vector(to_unsigned(character'pos(c), 7));
  end function;

begin

  process(clk)
    variable idx : integer;
  begin
    if rising_edge(clk) then
      idx := to_integer(unsigned(addr));
      if idx >= 0 and idx < ROM_SIZE then
        o_char <= char_to_slv(CHAR_ROM(idx));
      else
        o_char <= (others => '0');
      end if;
    end if;
  end process;

end rtl;
